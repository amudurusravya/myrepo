//------------------------------------------------------------------------------
// lookup table for square root unit
// this will have c0,c1 stored when x is [1 2) and 47:40 are used for table lookup
// sqrt_unit_lut_1.v
//
//------------------------------------------------------------------------------

module sqrt_unit_lut_1(
  input [5:0] addr,
  output [11:0] c1_sqrt1_out,
  output [19:0] c0_sqrt1_out
);

reg [11:0] c1_sqrt1;
reg [19:0] c0_sqrt1;

assign c0_sqrt1_out = c0_sqrt1;
assign c1_sqrt1_out = c1_sqrt1;

always @(addr) begin
  case(addr)
6'b000000 : c0_sqrt1 = 20'b00100000000111111100;
6'b000001 : c0_sqrt1 = 20'b00100000010111110011;
6'b000010 : c0_sqrt1 = 20'b00100000100111100100;
6'b000011 : c0_sqrt1 = 20'b00100000110111001101;
6'b000100 : c0_sqrt1 = 20'b00100001000110101111;
6'b000101 : c0_sqrt1 = 20'b00100001010110001000;
6'b000110 : c0_sqrt1 = 20'b00100001100101011101;
6'b000111 : c0_sqrt1 = 20'b00100001110100101001;
6'b001000 : c0_sqrt1 = 20'b00100010000011101110;
6'b001001 : c0_sqrt1 = 20'b00100010010010101101;
6'b001010 : c0_sqrt1 = 20'b00100010100001100101;
6'b001011 : c0_sqrt1 = 20'b00100010110000010111;
6'b001100 : c0_sqrt1 = 20'b00100010111111000010;
6'b001101 : c0_sqrt1 = 20'b00100011001101100111;
6'b001110 : c0_sqrt1 = 20'b00100011011100000111;
6'b001111 : c0_sqrt1 = 20'b00100011101010100010;
6'b010000 : c0_sqrt1 = 20'b00100011111000110101;
6'b010001 : c0_sqrt1 = 20'b00100100000111000101;
6'b010010 : c0_sqrt1 = 20'b00100100010101001101;
6'b010011 : c0_sqrt1 = 20'b00100100100011010001;
6'b010100 : c0_sqrt1 = 20'b00100100110001001110;
6'b010101 : c0_sqrt1 = 20'b00100100111111000111;
6'b010110 : c0_sqrt1 = 20'b00100101001100111011;
6'b010111 : c0_sqrt1 = 20'b00100101011010101001;
6'b011000 : c0_sqrt1 = 20'b00100101101000010010;
6'b011001 : c0_sqrt1 = 20'b00100101110101110101;
6'b011010 : c0_sqrt1 = 20'b00100110000011010100;
6'b011011 : c0_sqrt1 = 20'b00100110010000110000;
6'b011100 : c0_sqrt1 = 20'b00100110011110000110;
6'b011101 : c0_sqrt1 = 20'b00100110101011011000;
6'b011110 : c0_sqrt1 = 20'b00100110111000100100;
6'b011111 : c0_sqrt1 = 20'b00100111000101101101;
6'b100000 : c0_sqrt1 = 20'b00100111010010110001;
6'b100001 : c0_sqrt1 = 20'b00100111011111110000;
6'b100010 : c0_sqrt1 = 20'b00100111101100101101;
6'b100011 : c0_sqrt1 = 20'b00100111111001100100;
6'b100100 : c0_sqrt1 = 20'b00101000000110010110;
6'b100101 : c0_sqrt1 = 20'b00101000010011000101;
6'b100110 : c0_sqrt1 = 20'b00101000011111110010;
6'b100111 : c0_sqrt1 = 20'b00101000101100011001;
6'b101000 : c0_sqrt1 = 20'b00101000111000111011;
6'b101001 : c0_sqrt1 = 20'b00101001000101011011;
6'b101010 : c0_sqrt1 = 20'b00101001010001111000;
6'b101011 : c0_sqrt1 = 20'b00101001011110001111;
6'b101100 : c0_sqrt1 = 20'b00101001101010100100;
6'b101101 : c0_sqrt1 = 20'b00101001110110110100;
6'b101110 : c0_sqrt1 = 20'b00101010000011000001;
6'b101111 : c0_sqrt1 = 20'b00101010001111001001;
6'b110000 : c0_sqrt1 = 20'b00101010011011010001;
6'b110001 : c0_sqrt1 = 20'b00101010100111010100;
6'b110010 : c0_sqrt1 = 20'b00101010110011010010;
6'b110011 : c0_sqrt1 = 20'b00101010111111001111;
6'b110100 : c0_sqrt1 = 20'b00101011001011000111;
6'b110101 : c0_sqrt1 = 20'b00101011010110111101;
6'b110110 : c0_sqrt1 = 20'b00101011100010110000;
6'b110111 : c0_sqrt1 = 20'b00101011101110011110;
6'b111000 : c0_sqrt1 = 20'b00101011111010001001;
6'b111001 : c0_sqrt1 = 20'b00101100000101110001;
6'b111010 : c0_sqrt1 = 20'b00101100010001010111;
6'b111011 : c0_sqrt1 = 20'b00101100011100111010;
6'b111100 : c0_sqrt1 = 20'b00101100101000011011;
6'b111101 : c0_sqrt1 = 20'b00101100110011110110;
6'b111110 : c0_sqrt1 = 20'b00101100111111010010;
6'b111111 : c0_sqrt1 = 20'b00101101001010101000;
endcase
end
always @(addr) begin
  case(addr)
6'b000000 : c1_sqrt1 = 12'b000111111110;
6'b000001 : c1_sqrt1 = 12'b000111111010;
6'b000010 : c1_sqrt1 = 12'b000111110110;
6'b000011 : c1_sqrt1 = 12'b000111110010;
6'b000100 : c1_sqrt1 = 12'b000111101110;
6'b000101 : c1_sqrt1 = 12'b000111101011;
6'b000110 : c1_sqrt1 = 12'b000111100111;
6'b000111 : c1_sqrt1 = 12'b000111100100;
6'b001000 : c1_sqrt1 = 12'b000111100001;
6'b001001 : c1_sqrt1 = 12'b000111011101;
6'b001010 : c1_sqrt1 = 12'b000111011010;
6'b001011 : c1_sqrt1 = 12'b000111010111;
6'b001100 : c1_sqrt1 = 12'b000111010100;
6'b001101 : c1_sqrt1 = 12'b000111010001;
6'b001110 : c1_sqrt1 = 12'b000111001110;
6'b001111 : c1_sqrt1 = 12'b000111001011;
6'b010000 : c1_sqrt1 = 12'b000111001000;
6'b010001 : c1_sqrt1 = 12'b000111000101;
6'b010010 : c1_sqrt1 = 12'b000111000010;
6'b010011 : c1_sqrt1 = 12'b000111000000;
6'b010100 : c1_sqrt1 = 12'b000110111101;
6'b010101 : c1_sqrt1 = 12'b000110111010;
6'b010110 : c1_sqrt1 = 12'b000110111000;
6'b010111 : c1_sqrt1 = 12'b000110110101;
6'b011000 : c1_sqrt1 = 12'b000110110011;
6'b011001 : c1_sqrt1 = 12'b000110110000;
6'b011010 : c1_sqrt1 = 12'b000110101110;
6'b011011 : c1_sqrt1 = 12'b000110101100;
6'b011100 : c1_sqrt1 = 12'b000110101001;
6'b011101 : c1_sqrt1 = 12'b000110100111;
6'b011110 : c1_sqrt1 = 12'b000110100101;
6'b011111 : c1_sqrt1 = 12'b000110100011;
6'b100000 : c1_sqrt1 = 12'b000110100000;
6'b100001 : c1_sqrt1 = 12'b000110011110;
6'b100010 : c1_sqrt1 = 12'b000110011100;
6'b100011 : c1_sqrt1 = 12'b000110011010;
6'b100100 : c1_sqrt1 = 12'b000110011000;
6'b100101 : c1_sqrt1 = 12'b000110010110;
6'b100110 : c1_sqrt1 = 12'b000110010100;
6'b100111 : c1_sqrt1 = 12'b000110010010;
6'b101000 : c1_sqrt1 = 12'b000110010000;
6'b101001 : c1_sqrt1 = 12'b000110001110;
6'b101010 : c1_sqrt1 = 12'b000110001100;
6'b101011 : c1_sqrt1 = 12'b000110001011;
6'b101100 : c1_sqrt1 = 12'b000110001001;
6'b101101 : c1_sqrt1 = 12'b000110000111;
6'b101110 : c1_sqrt1 = 12'b000110000101;
6'b101111 : c1_sqrt1 = 12'b000110000011;
6'b110000 : c1_sqrt1 = 12'b000110000010;
6'b110001 : c1_sqrt1 = 12'b000110000000;
6'b110010 : c1_sqrt1 = 12'b000101111110;
6'b110011 : c1_sqrt1 = 12'b000101111101;
6'b110100 : c1_sqrt1 = 12'b000101111011;
6'b110101 : c1_sqrt1 = 12'b000101111001;
6'b110110 : c1_sqrt1 = 12'b000101111000;
6'b110111 : c1_sqrt1 = 12'b000101110110;
6'b111000 : c1_sqrt1 = 12'b000101110101;
6'b111001 : c1_sqrt1 = 12'b000101110011;
6'b111010 : c1_sqrt1 = 12'b000101110010;
6'b111011 : c1_sqrt1 = 12'b000101110000;
6'b111100 : c1_sqrt1 = 12'b000101101111;
6'b111101 : c1_sqrt1 = 12'b000101101101;
6'b111110 : c1_sqrt1 = 12'b000101101100;
6'b111111 : c1_sqrt1 = 12'b000101101010;
endcase
end
endmodule
