//------------------------------------------------------------------------------
// lookup table for logarithm unit
// this will have c0,c1,c2 stored and 47:40 are used for table lookup
// log_unit_lut.v
//
//------------------------------------------------------------------------------

module log_unit_lut(
  input [7:0] addr,
  output [12:0] c2_log_out,
  output [21:0] c1_log_out,
  output [29:0] c0_log_out
);

reg [12:0] c2_log;
reg [21:0] c1_log;
reg [29:0] c0_log;

assign c0_log_out = c0_log;
assign c1_log_out = c1_log;
assign c2_log_out = c2_log;

always @(addr) begin
  case(addr)
8'b00000000 : c2_log = 0001111111100;
8'b00000001 : c2_log = 0001111110100;
8'b00000010 : c2_log = 0001111101100;
8'b00000011 : c2_log = 0001111100100;
8'b00000100 : c2_log = 0001111011100;
8'b00000101 : c2_log = 0001111010101;
8'b00000110 : c2_log = 0001111001101;
8'b00000111 : c2_log = 0001111000110;
8'b00001000 : c2_log = 0001110111111;
8'b00001001 : c2_log = 0001110111000;
8'b00001010 : c2_log = 0001110110000;
8'b00001011 : c2_log = 0001110101001;
8'b00001100 : c2_log = 0001110100010;
8'b00001101 : c2_log = 0001110011011;
8'b00001110 : c2_log = 0001110010101;
8'b00001111 : c2_log = 0001110001110;
8'b00010000 : c2_log = 0001110000111;
8'b00010001 : c2_log = 0001110000001;
8'b00010010 : c2_log = 0001101111010;
8'b00010011 : c2_log = 0001101110100;
8'b00010100 : c2_log = 0001101101101;
8'b00010101 : c2_log = 0001101100111;
8'b00010110 : c2_log = 0001101100001;
8'b00010111 : c2_log = 0001101011011;
8'b00011000 : c2_log = 0001101010100;
8'b00011001 : c2_log = 0001101001110;
8'b00011010 : c2_log = 0001101001000;
8'b00011011 : c2_log = 0001101000010;
8'b00011100 : c2_log = 0001100111101;
8'b00011101 : c2_log = 0001100110111;
8'b00011110 : c2_log = 0001100110001;
8'b00011111 : c2_log = 0001100101011;
8'b00100000 : c2_log = 0001100100110;
8'b00100001 : c2_log = 0001100100000;
8'b00100010 : c2_log = 0001100011011;
8'b00100011 : c2_log = 0001100010101;
8'b00100100 : c2_log = 0001100010000;
8'b00100101 : c2_log = 0001100001011;
8'b00100110 : c2_log = 0001100000101;
8'b00100111 : c2_log = 0001100000000;
8'b00101000 : c2_log = 0001011111011;
8'b00101001 : c2_log = 0001011110110;
8'b00101010 : c2_log = 0001011110001;
8'b00101011 : c2_log = 0001011101100;
8'b00101100 : c2_log = 0001011100111;
8'b00101101 : c2_log = 0001011100010;
8'b00101110 : c2_log = 0001011011101;
8'b00101111 : c2_log = 0001011011000;
8'b00110000 : c2_log = 0001011010011;
8'b00110001 : c2_log = 0001011001111;
8'b00110010 : c2_log = 0001011001010;
8'b00110011 : c2_log = 0001011000101;
8'b00110100 : c2_log = 0001011000001;
8'b00110101 : c2_log = 0001010111100;
8'b00110110 : c2_log = 0001010111000;
8'b00110111 : c2_log = 0001010110011;
8'b00111000 : c2_log = 0001010101111;
8'b00111001 : c2_log = 0001010101010;
8'b00111010 : c2_log = 0001010100110;
8'b00111011 : c2_log = 0001010100010;
8'b00111100 : c2_log = 0001010011101;
8'b00111101 : c2_log = 0001010011001;
8'b00111110 : c2_log = 0001010010101;
8'b00111111 : c2_log = 0001010010001;
8'b01000000 : c2_log = 0001010001101;
8'b01000001 : c2_log = 0001010001001;
8'b01000010 : c2_log = 0001010000101;
8'b01000011 : c2_log = 0001010000001;
8'b01000100 : c2_log = 0001001111101;
8'b01000101 : c2_log = 0001001111001;
8'b01000110 : c2_log = 0001001110101;
8'b01000111 : c2_log = 0001001110001;
8'b01001000 : c2_log = 0001001101101;
8'b01001001 : c2_log = 0001001101010;
8'b01001010 : c2_log = 0001001100110;
8'b01001011 : c2_log = 0001001100010;
8'b01001100 : c2_log = 0001001011111;
8'b01001101 : c2_log = 0001001011011;
8'b01001110 : c2_log = 0001001010111;
8'b01001111 : c2_log = 0001001010100;
8'b01010000 : c2_log = 0001001010000;
8'b01010001 : c2_log = 0001001001101;
8'b01010010 : c2_log = 0001001001001;
8'b01010011 : c2_log = 0001001000110;
8'b01010100 : c2_log = 0001001000010;
8'b01010101 : c2_log = 0001000111111;
8'b01010110 : c2_log = 0001000111100;
8'b01010111 : c2_log = 0001000111000;
8'b01011000 : c2_log = 0001000110101;
8'b01011001 : c2_log = 0001000110010;
8'b01011010 : c2_log = 0001000101110;
8'b01011011 : c2_log = 0001000101011;
8'b01011100 : c2_log = 0001000101000;
8'b01011101 : c2_log = 0001000100101;
8'b01011110 : c2_log = 0001000100010;
8'b01011111 : c2_log = 0001000011111;
8'b01100000 : c2_log = 0001000011100;
8'b01100001 : c2_log = 0001000011001;
8'b01100010 : c2_log = 0001000010110;
8'b01100011 : c2_log = 0001000010011;
8'b01100100 : c2_log = 0001000010000;
8'b01100101 : c2_log = 0001000001101;
8'b01100110 : c2_log = 0001000001010;
8'b01100111 : c2_log = 0001000000111;
8'b01101000 : c2_log = 0001000000100;
8'b01101001 : c2_log = 0001000000001;
8'b01101010 : c2_log = 0000111111110;
8'b01101011 : c2_log = 0000111111011;
8'b01101100 : c2_log = 0000111111001;
8'b01101101 : c2_log = 0000111110110;
8'b01101110 : c2_log = 0000111110011;
8'b01101111 : c2_log = 0000111110000;
8'b01110000 : c2_log = 0000111101110;
8'b01110001 : c2_log = 0000111101011;
8'b01110010 : c2_log = 0000111101000;
8'b01110011 : c2_log = 0000111100110;
8'b01110100 : c2_log = 0000111100011;
8'b01110101 : c2_log = 0000111100001;
8'b01110110 : c2_log = 0000111011110;
8'b01110111 : c2_log = 0000111011011;
8'b01111000 : c2_log = 0000111011001;
8'b01111001 : c2_log = 0000111010110;
8'b01111010 : c2_log = 0000111010100;
8'b01111011 : c2_log = 0000111010001;
8'b01111100 : c2_log = 0000111001111;
8'b01111101 : c2_log = 0000111001101;
8'b01111110 : c2_log = 0000111001010;
8'b01111111 : c2_log = 0000111001000;
8'b10000000 : c2_log = 0000111000101;
8'b10000001 : c2_log = 0000111000011;
8'b10000010 : c2_log = 0000111000001;
8'b10000011 : c2_log = 0000110111110;
8'b10000100 : c2_log = 0000110111100;
8'b10000101 : c2_log = 0000110111010;
8'b10000110 : c2_log = 0000110111000;
8'b10000111 : c2_log = 0000110110101;
8'b10001000 : c2_log = 0000110110011;
8'b10001001 : c2_log = 0000110110001;
8'b10001010 : c2_log = 0000110101111;
8'b10001011 : c2_log = 0000110101101;
8'b10001100 : c2_log = 0000110101010;
8'b10001101 : c2_log = 0000110101000;
8'b10001110 : c2_log = 0000110100110;
8'b10001111 : c2_log = 0000110100100;
8'b10010000 : c2_log = 0000110100010;
8'b10010001 : c2_log = 0000110100000;
8'b10010010 : c2_log = 0000110011110;
8'b10010011 : c2_log = 0000110011100;
8'b10010100 : c2_log = 0000110011010;
8'b10010101 : c2_log = 0000110011000;
8'b10010110 : c2_log = 0000110010110;
8'b10010111 : c2_log = 0000110010100;
8'b10011000 : c2_log = 0000110010010;
8'b10011001 : c2_log = 0000110010000;
8'b10011010 : c2_log = 0000110001110;
8'b10011011 : c2_log = 0000110001100;
8'b10011100 : c2_log = 0000110001010;
8'b10011101 : c2_log = 0000110001000;
8'b10011110 : c2_log = 0000110000110;
8'b10011111 : c2_log = 0000110000100;
8'b10100000 : c2_log = 0000110000010;
8'b10100001 : c2_log = 0000110000001;
8'b10100010 : c2_log = 0000101111111;
8'b10100011 : c2_log = 0000101111101;
8'b10100100 : c2_log = 0000101111011;
8'b10100101 : c2_log = 0000101111001;
8'b10100110 : c2_log = 0000101110111;
8'b10100111 : c2_log = 0000101110110;
8'b10101000 : c2_log = 0000101110100;
8'b10101001 : c2_log = 0000101110010;
8'b10101010 : c2_log = 0000101110000;
8'b10101011 : c2_log = 0000101101111;
8'b10101100 : c2_log = 0000101101101;
8'b10101101 : c2_log = 0000101101011;
8'b10101110 : c2_log = 0000101101010;
8'b10101111 : c2_log = 0000101101000;
8'b10110000 : c2_log = 0000101100110;
8'b10110001 : c2_log = 0000101100101;
8'b10110010 : c2_log = 0000101100011;
8'b10110011 : c2_log = 0000101100001;
8'b10110100 : c2_log = 0000101100000;
8'b10110101 : c2_log = 0000101011110;
8'b10110110 : c2_log = 0000101011101;
8'b10110111 : c2_log = 0000101011011;
8'b10111000 : c2_log = 0000101011001;
8'b10111001 : c2_log = 0000101011000;
8'b10111010 : c2_log = 0000101010110;
8'b10111011 : c2_log = 0000101010101;
8'b10111100 : c2_log = 0000101010011;
8'b10111101 : c2_log = 0000101010010;
8'b10111110 : c2_log = 0000101010000;
8'b10111111 : c2_log = 0000101001111;
8'b11000000 : c2_log = 0000101001101;
8'b11000001 : c2_log = 0000101001100;
8'b11000010 : c2_log = 0000101001010;
8'b11000011 : c2_log = 0000101001001;
8'b11000100 : c2_log = 0000101000111;
8'b11000101 : c2_log = 0000101000110;
8'b11000110 : c2_log = 0000101000100;
8'b11000111 : c2_log = 0000101000011;
8'b11001000 : c2_log = 0000101000010;
8'b11001001 : c2_log = 0000101000000;
8'b11001010 : c2_log = 0000100111111;
8'b11001011 : c2_log = 0000100111101;
8'b11001100 : c2_log = 0000100111100;
8'b11001101 : c2_log = 0000100111011;
8'b11001110 : c2_log = 0000100111001;
8'b11001111 : c2_log = 0000100111000;
8'b11010000 : c2_log = 0000100110111;
8'b11010001 : c2_log = 0000100110101;
8'b11010010 : c2_log = 0000100110100;
8'b11010011 : c2_log = 0000100110011;
8'b11010100 : c2_log = 0000100110001;
8'b11010101 : c2_log = 0000100110000;
8'b11010110 : c2_log = 0000100101111;
8'b11010111 : c2_log = 0000100101101;
8'b11011000 : c2_log = 0000100101100;
8'b11011001 : c2_log = 0000100101011;
8'b11011010 : c2_log = 0000100101010;
8'b11011011 : c2_log = 0000100101000;
8'b11011100 : c2_log = 0000100100111;
8'b11011101 : c2_log = 0000100100110;
8'b11011110 : c2_log = 0000100100101;
8'b11011111 : c2_log = 0000100100011;
8'b11100000 : c2_log = 0000100100010;
8'b11100001 : c2_log = 0000100100001;
8'b11100010 : c2_log = 0000100100000;
8'b11100011 : c2_log = 0000100011111;
8'b11100100 : c2_log = 0000100011101;
8'b11100101 : c2_log = 0000100011100;
8'b11100110 : c2_log = 0000100011011;
8'b11100111 : c2_log = 0000100011010;
8'b11101000 : c2_log = 0000100011001;
8'b11101001 : c2_log = 0000100011000;
8'b11101010 : c2_log = 0000100010110;
8'b11101011 : c2_log = 0000100010101;
8'b11101100 : c2_log = 0000100010100;
8'b11101101 : c2_log = 0000100010011;
8'b11101110 : c2_log = 0000100010010;
8'b11101111 : c2_log = 0000100010001;
8'b11110000 : c2_log = 0000100010000;
8'b11110001 : c2_log = 0000100001111;
8'b11110010 : c2_log = 0000100001110;
8'b11110011 : c2_log = 0000100001100;
8'b11110100 : c2_log = 0000100001011;
8'b11110101 : c2_log = 0000100001010;
8'b11110110 : c2_log = 0000100001001;
8'b11110111 : c2_log = 0000100001000;
8'b11111000 : c2_log = 0000100000111;
8'b11111001 : c2_log = 0000100000110;
8'b11111010 : c2_log = 0000100000101;
8'b11111011 : c2_log = 0000100000100;
8'b11111100 : c2_log = 0000100000011;
8'b11111101 : c2_log = 0000100000010;
8'b11111110 : c2_log = 0000100000001;
8'b11111111 : c2_log = 0000100000000;
endcase
end

always @(addr) begin
  case(addr)
8'b00000000 : c1_log = 22'b1111111111000000000110;
8'b00000001 : c1_log = 22'b1111111101000001111100;
8'b00000010 : c1_log = 22'b1111111011000011110010;
8'b00000011 : c1_log = 22'b1111111001000101101000;
8'b00000100 : c1_log = 22'b1111110111001010110000;
8'b00000101 : c1_log = 22'b1111110101001110001110;
8'b00000110 : c1_log = 22'b1111110011010100111111;
8'b00000111 : c1_log = 22'b1111110001011011110000;
8'b00001000 : c1_log = 22'b1111101111100010100000;
8'b00001001 : c1_log = 22'b1111101101101010111001;
8'b00001010 : c1_log = 22'b1111101011110100111100;
8'b00001011 : c1_log = 22'b1111101001111110111110;
8'b00001100 : c1_log = 22'b1111101000001010101001;
8'b00001101 : c1_log = 22'b1111100110010110010100;
8'b00001110 : c1_log = 22'b1111100100100011101000;
8'b00001111 : c1_log = 22'b1111100010110000111100;
8'b00010000 : c1_log = 22'b1111100000111111111001;
8'b00010001 : c1_log = 22'b1111011111001110110110;
8'b00010010 : c1_log = 22'b1111011101011111011011;
8'b00010011 : c1_log = 22'b1111011011110000000001;
8'b00010100 : c1_log = 22'b1111011010000010010000;
8'b00010101 : c1_log = 22'b1111011000010100011110;
8'b00010110 : c1_log = 22'b1111010110101000010110;
8'b00010111 : c1_log = 22'b1111010100111100001101;
8'b00011000 : c1_log = 22'b1111010011010001101101;
8'b00011001 : c1_log = 22'b1111010001100111001110;
8'b00011010 : c1_log = 22'b1111001111111110010111;
8'b00011011 : c1_log = 22'b1111001110010101100000;
8'b00011100 : c1_log = 22'b1111001100101110010010;
8'b00011101 : c1_log = 22'b1111001011000101011011;
8'b00011110 : c1_log = 22'b1111001001011111110110;
8'b00011111 : c1_log = 22'b1111000111111010010000;
8'b00100000 : c1_log = 22'b1111000110010100101011;
8'b00100001 : c1_log = 22'b1111000100110000101111;
8'b00100010 : c1_log = 22'b1111000011001100110011;
8'b00100011 : c1_log = 22'b1111000001101000110110;
8'b00100100 : c1_log = 22'b1111000000000110100011;
8'b00100101 : c1_log = 22'b1110111110100101111000;
8'b00100110 : c1_log = 22'b1110111101000011100101;
8'b00100111 : c1_log = 22'b1110111011100100100011;
8'b00101000 : c1_log = 22'b1110111010000011111001;
8'b00101001 : c1_log = 22'b1110111000100100110111;
8'b00101010 : c1_log = 22'b1110110111000101110101;
8'b00101011 : c1_log = 22'b1110110101101000011100;
8'b00101100 : c1_log = 22'b1110110100001011000011;
8'b00101101 : c1_log = 22'b1110110010101111010011;
8'b00101110 : c1_log = 22'b1110110001010011100011;
8'b00101111 : c1_log = 22'b1110101111110111110011;
8'b00110000 : c1_log = 22'b1110101110011100000011;
8'b00110001 : c1_log = 22'b1110101101000001111100;
8'b00110010 : c1_log = 22'b1110101011101001011110;
8'b00110011 : c1_log = 22'b1110101010001111010111;
8'b00110100 : c1_log = 22'b1110101000110110111000;
8'b00110101 : c1_log = 22'b1110100111100000000011;
8'b00110110 : c1_log = 22'b1110100110001001001101;
8'b00110111 : c1_log = 22'b1110100100110010011000;
8'b00111000 : c1_log = 22'b1110100011011011100010;
8'b00111001 : c1_log = 22'b1110100010000110010110;
8'b00111010 : c1_log = 22'b1110100000110001001001;
8'b00111011 : c1_log = 22'b1110011111011011111101;
8'b00111100 : c1_log = 22'b1110011110001000011001;
8'b00111101 : c1_log = 22'b1110011100110100110101;
8'b00111110 : c1_log = 22'b1110011011100001010001;
8'b00111111 : c1_log = 22'b1110011010001111010111;
8'b01000000 : c1_log = 22'b1110011000111101011100;
8'b01000001 : c1_log = 22'b1110010111101011100001;
8'b01000010 : c1_log = 22'b1110010110011011001111;
8'b01000011 : c1_log = 22'b1110010101001010111101;
8'b01000100 : c1_log = 22'b1110010011111010101011;
8'b01000101 : c1_log = 22'b1110010010101100000010;
8'b01000110 : c1_log = 22'b1110010001011011110000;
8'b01000111 : c1_log = 22'b1110010000001110101111;
8'b01001000 : c1_log = 22'b1110001111000000000110;
8'b01001001 : c1_log = 22'b1110001101110011000110;
8'b01001010 : c1_log = 22'b1110001100100110000101;
8'b01001011 : c1_log = 22'b1110001011011001000101;
8'b01001100 : c1_log = 22'b1110001010001101101110;
8'b01001101 : c1_log = 22'b1110001001000000101101;
8'b01001110 : c1_log = 22'b1110000111110101010110;
8'b01001111 : c1_log = 22'b1110000110101011100111;
8'b01010000 : c1_log = 22'b1110000101100000010000;
8'b01010001 : c1_log = 22'b1110000100010110100001;
8'b01010010 : c1_log = 22'b1110000011001110011100;
8'b01010011 : c1_log = 22'b1110000010000100101101;
8'b01010100 : c1_log = 22'b1110000000111100100111;
8'b01010101 : c1_log = 22'b1101111111110100100001;
8'b01010110 : c1_log = 22'b1101111110101100011100;
8'b01010111 : c1_log = 22'b1101111101100100010110;
8'b01011000 : c1_log = 22'b1101111100011101111001;
8'b01011001 : c1_log = 22'b1101111011010111011100;
8'b01011010 : c1_log = 22'b1101111010010000111111;
8'b01011011 : c1_log = 22'b1101111001001100001011;
8'b01011100 : c1_log = 22'b1101111000000111010111;
8'b01011101 : c1_log = 22'b1101110111000010100011;
8'b01011110 : c1_log = 22'b1101110101111101101111;
8'b01011111 : c1_log = 22'b1101110100111000111011;
8'b01100000 : c1_log = 22'b1101110011110101110000;
8'b01100001 : c1_log = 22'b1101110010110010100101;
8'b01100010 : c1_log = 22'b1101110001101111011010;
8'b01100011 : c1_log = 22'b1101110000101100001111;
8'b01100100 : c1_log = 22'b1101101111101010101100;
8'b01100101 : c1_log = 22'b1101101110101001001010;
8'b01100110 : c1_log = 22'b1101101101100111101000;
8'b01100111 : c1_log = 22'b1101101100100110000101;
8'b01101000 : c1_log = 22'b1101101011100110001100;
8'b01101001 : c1_log = 22'b1101101010100100101010;
8'b01101010 : c1_log = 22'b1101101001100100110000;
8'b01101011 : c1_log = 22'b1101101000100100110111;
8'b01101100 : c1_log = 22'b1101100111100110100110;
8'b01101101 : c1_log = 22'b1101100110100110101101;
8'b01101110 : c1_log = 22'b1101100101101000011100;
8'b01101111 : c1_log = 22'b1101100100101010001100;
8'b01110000 : c1_log = 22'b1101100011101011111011;
8'b01110001 : c1_log = 22'b1101100010101111010011;
8'b01110010 : c1_log = 22'b1101100001110001000011;
8'b01110011 : c1_log = 22'b1101100000110100011011;
8'b01110100 : c1_log = 22'b1101011111110111110011;
8'b01110101 : c1_log = 22'b1101011110111011001011;
8'b01110110 : c1_log = 22'b1101011110000000001101;
8'b01110111 : c1_log = 22'b1101011101000011100101;
8'b01111000 : c1_log = 22'b1101011100001000100110;
8'b01111001 : c1_log = 22'b1101011011001101100111;
8'b01111010 : c1_log = 22'b1101011010010010101000;
8'b01111011 : c1_log = 22'b1101011001010111101001;
8'b01111100 : c1_log = 22'b1101011000011110010011;
8'b01111101 : c1_log = 22'b1101010111100100111101;
8'b01111110 : c1_log = 22'b1101010110101011100111;
8'b01111111 : c1_log = 22'b1101010101110010010001;
8'b10000000 : c1_log = 22'b1101010100111000111011;
8'b10000001 : c1_log = 22'b1101010011111111100101;
8'b10000010 : c1_log = 22'b1101010011000111111000;
8'b10000011 : c1_log = 22'b1101010010010000001011;
8'b10000100 : c1_log = 22'b1101010001011000011110;
8'b10000101 : c1_log = 22'b1101010000100000110001;
8'b10000110 : c1_log = 22'b1101001111101001000011;
8'b10000111 : c1_log = 22'b1101001110110010111111;
8'b10001000 : c1_log = 22'b1101001101111100111011;
8'b10001001 : c1_log = 22'b1101001101000101001110;
8'b10001010 : c1_log = 22'b1101001100001111001001;
8'b10001011 : c1_log = 22'b1101001011011010101110;
8'b10001100 : c1_log = 22'b1101001010100100101010;
8'b10001101 : c1_log = 22'b1101001001110000001110;
8'b10001110 : c1_log = 22'b1101001000111010001010;
8'b10001111 : c1_log = 22'b1101001000000101101111;
8'b10010000 : c1_log = 22'b1101000111010001010011;
8'b10010001 : c1_log = 22'b1101000110011100111000;
8'b10010010 : c1_log = 22'b1101000101101010000101;
8'b10010011 : c1_log = 22'b1101000100110101101010;
8'b10010100 : c1_log = 22'b1101000100000010110111;
8'b10010101 : c1_log = 22'b1101000011001110011100;
8'b10010110 : c1_log = 22'b1101000010011011101001;
8'b10010111 : c1_log = 22'b1101000001101000110110;
8'b10011000 : c1_log = 22'b1101000000110111101101;
8'b10011001 : c1_log = 22'b1101000000000100111010;
8'b10011010 : c1_log = 22'b1100111111010011110000;
8'b10011011 : c1_log = 22'b1100111110100000111110;
8'b10011100 : c1_log = 22'b1100111101101111110100;
8'b10011101 : c1_log = 22'b1100111100111110101010;
8'b10011110 : c1_log = 22'b1100111100001101100001;
8'b10011111 : c1_log = 22'b1100111011011110000000;
8'b10100000 : c1_log = 22'b1100111010101100110110;
8'b10100001 : c1_log = 22'b1100111001111011101100;
8'b10100010 : c1_log = 22'b1100111001001100001011;
8'b10100011 : c1_log = 22'b1100111000011100101011;
8'b10100100 : c1_log = 22'b1100110111101101001010;
8'b10100101 : c1_log = 22'b1100110110111101101001;
8'b10100110 : c1_log = 22'b1100110110001110001000;
8'b10100111 : c1_log = 22'b1100110101100000010000;
8'b10101000 : c1_log = 22'b1100110100110000101111;
8'b10101001 : c1_log = 22'b1100110100000010110111;
8'b10101010 : c1_log = 22'b1100110011010100111111;
8'b10101011 : c1_log = 22'b1100110010100111000111;
8'b10101100 : c1_log = 22'b1100110001111001001111;
8'b10101101 : c1_log = 22'b1100110001001011010111;
8'b10101110 : c1_log = 22'b1100110000011101011111;
8'b10101111 : c1_log = 22'b1100101111110001010000;
8'b10110000 : c1_log = 22'b1100101111000011011000;
8'b10110001 : c1_log = 22'b1100101110010111001001;
8'b10110010 : c1_log = 22'b1100101101101010111001;
8'b10110011 : c1_log = 22'b1100101100111110101010;
8'b10110100 : c1_log = 22'b1100101100010010011011;
8'b10110101 : c1_log = 22'b1100101011100110001100;
8'b10110110 : c1_log = 22'b1100101010111001111101;
8'b10110111 : c1_log = 22'b1100101010001111010111;
8'b10111000 : c1_log = 22'b1100101001100011000111;
8'b10111001 : c1_log = 22'b1100101000111000100001;
8'b10111010 : c1_log = 22'b1100101000001101111011;
8'b10111011 : c1_log = 22'b1100100111100011010100;
8'b10111100 : c1_log = 22'b1100100110111000101110;
8'b10111101 : c1_log = 22'b1100100110001110001000;
8'b10111110 : c1_log = 22'b1100100101100011100010;
8'b10111111 : c1_log = 22'b1100100100111000111011;
8'b11000000 : c1_log = 22'b1100100100001111111110;
8'b11000001 : c1_log = 22'b1100100011100101011000;
8'b11000010 : c1_log = 22'b1100100010111100011010;
8'b11000011 : c1_log = 22'b1100100010010011011101;
8'b11000100 : c1_log = 22'b1100100001101010011111;
8'b11000101 : c1_log = 22'b1100100001000001100010;
8'b11000110 : c1_log = 22'b1100100000011000100100;
8'b11000111 : c1_log = 22'b1100011111101111100111;
8'b11001000 : c1_log = 22'b1100011111001000010010;
8'b11001001 : c1_log = 22'b1100011110011111010101;
8'b11001010 : c1_log = 22'b1100011101111000000000;
8'b11001011 : c1_log = 22'b1100011101010000101100;
8'b11001100 : c1_log = 22'b1100011100100111101110;
8'b11001101 : c1_log = 22'b1100011100000000011010;
8'b11001110 : c1_log = 22'b1100011011011001000101;
8'b11001111 : c1_log = 22'b1100011010110001110001;
8'b11010000 : c1_log = 22'b1100011010001100000101;
8'b11010001 : c1_log = 22'b1100011001100100110000;
8'b11010010 : c1_log = 22'b1100011000111101011100;
8'b11010011 : c1_log = 22'b1100011000010111110000;
8'b11010100 : c1_log = 22'b1100010111110010000100;
8'b11010101 : c1_log = 22'b1100010111001010110000;
8'b11010110 : c1_log = 22'b1100010110100101000100;
8'b11010111 : c1_log = 22'b1100010101111111011000;
8'b11011000 : c1_log = 22'b1100010101011001101100;
8'b11011001 : c1_log = 22'b1100010100110100000001;
8'b11011010 : c1_log = 22'b1100010100001110010101;
8'b11011011 : c1_log = 22'b1100010011101010010010;
8'b11011100 : c1_log = 22'b1100010011000100100110;
8'b11011101 : c1_log = 22'b1100010010100000100100;
8'b11011110 : c1_log = 22'b1100010001111010111000;
8'b11011111 : c1_log = 22'b1100010001010110110101;
8'b11100000 : c1_log = 22'b1100010000110010110010;
8'b11100001 : c1_log = 22'b1100010000001101000110;
8'b11100010 : c1_log = 22'b1100001111101001000011;
8'b11100011 : c1_log = 22'b1100001111000101000001;
8'b11100100 : c1_log = 22'b1100001110100010100111;
8'b11100101 : c1_log = 22'b1100001101111110100100;
8'b11100110 : c1_log = 22'b1100001101011010100001;
8'b11100111 : c1_log = 22'b1100001100111000000111;
8'b11101000 : c1_log = 22'b1100001100010100000100;
8'b11101001 : c1_log = 22'b1100001011110001101010;
8'b11101010 : c1_log = 22'b1100001011001101100111;
8'b11101011 : c1_log = 22'b1100001010101011001101;
8'b11101100 : c1_log = 22'b1100001010001000110011;
8'b11101101 : c1_log = 22'b1100001001100110011001;
8'b11101110 : c1_log = 22'b1100001001000011111111;
8'b11101111 : c1_log = 22'b1100001000100001100101;
8'b11110000 : c1_log = 22'b1100000111111111001011;
8'b11110001 : c1_log = 22'b1100000111011100110001;
8'b11110010 : c1_log = 22'b1100000110111100000000;
8'b11110011 : c1_log = 22'b1100000110011001100110;
8'b11110100 : c1_log = 22'b1100000101111000110101;
8'b11110101 : c1_log = 22'b1100000101010110011011;
8'b11110110 : c1_log = 22'b1100000100110101101010;
8'b11110111 : c1_log = 22'b1100000100010100111000;
8'b11111000 : c1_log = 22'b1100000011110100000111;
8'b11111001 : c1_log = 22'b1100000011010011010110;
8'b11111010 : c1_log = 22'b1100000010110010100101;
8'b11111011 : c1_log = 22'b1100000010010001110100;
8'b11111100 : c1_log = 22'b1100000001110001000011;
8'b11111101 : c1_log = 22'b1100000001010000010010;
8'b11111110 : c1_log = 22'b1100000000101111100000;
8'b11111111 : c1_log = 22'b1100000000010000011000;
endcase
end
always @(addr) begin
  case(addr)
8'b00000000 : c0_log = 30'b010111111110000011011110110100;
8'b00000001 : c0_log = 30'b010111111010000011111001000010;
8'b00000010 : c0_log = 30'b010111110110000100010011010000;
8'b00000011 : c0_log = 30'b010111110010000100101101011101;
8'b00000100 : c0_log = 30'b010111101110001011101011000111;
8'b00000101 : c0_log = 30'b010111101010001100000101010100;
8'b00000110 : c0_log = 30'b010111100110010011000010111110;
8'b00000111 : c0_log = 30'b010111100010011010000000100111;
8'b00001000 : c0_log = 30'b010111011110100000111110010000;
8'b00001001 : c0_log = 30'b010111011010101110011111010101;
8'b00001010 : c0_log = 30'b010111010110110101011100111110;
8'b00001011 : c0_log = 30'b010111010011000010111110000011;
8'b00001100 : c0_log = 30'b010111001111001001111011101100;
8'b00001101 : c0_log = 30'b010111001011010111011100110001;
8'b00001110 : c0_log = 30'b010111000111100100111101110110;
8'b00001111 : c0_log = 30'b010111000011110010011110111011;
8'b00010000 : c0_log = 30'b010111                        ;
8'b00010001 : c0_log = 30'b010110111100010100000100100000;
8'b00010010 : c0_log = 30'b010110111000100001100101100101;
8'b00010011 : c0_log = 30'b010110110100110101101010000101;
8'b00010100 : c0_log = 30'b010110110001001001101110100101;
8'b00010101 : c0_log = 30'b010110101101011101110011000110;
8'b00010110 : c0_log = 30'b010110101001110001110111100110;
8'b00010111 : c0_log = 30'b010110100110000101111100000110;
8'b00011000 : c0_log = 30'b010110100010011010000000100111;
8'b00011001 : c0_log = 30'b010110011110101110000101000111;
8'b00011010 : c0_log = 30'b010110011011001000101101000011;
8'b00011011 : c0_log = 30'b010110010111100011010100111111;
8'b00011100 : c0_log = 30'b010110010011110111011001011111;
8'b00011101 : c0_log = 30'b010110010000010010000001011011;
8'b00011110 : c0_log = 30'b010110001100101100101001010111;
8'b00011111 : c0_log = 30'b010110001001001101110100101111;
8'b00100000 : c0_log = 30'b010110000101101000011100101011;
8'b00100001 : c0_log = 30'b010110000010000011000100100110;
8'b00100010 : c0_log = 30'b010101111110100100001111111110;
8'b00100011 : c0_log = 30'b010101111010111110110111111010;
8'b00100100 : c0_log = 30'b010101110111100000000011010001;
8'b00100101 : c0_log = 30'b010101110100000001001110101001;
8'b00100110 : c0_log = 30'b010101110000100010011010000000;
8'b00100111 : c0_log = 30'b010101101101000011100101011000;
8'b00101000 : c0_log = 30'b010101101001100100110000101111;
8'b00101001 : c0_log = 30'b010101100110001100011111100010;
8'b00101010 : c0_log = 30'b010101100010101101101010111001;
8'b00101011 : c0_log = 30'b010101011111010101011001101100;
8'b00101100 : c0_log = 30'b010101011011110110100101000100;
8'b00101101 : c0_log = 30'b010101011000011110010011110111;
8'b00101110 : c0_log = 30'b010101010101000110000010101010;
8'b00101111 : c0_log = 30'b010101010001101101110001011101;
8'b00110000 : c0_log = 30'b010101001110010101100000010000;
8'b00110001 : c0_log = 30'b010101001010111101001111000011;
8'b00110010 : c0_log = 30'b010101000111101011100001010001;
8'b00110011 : c0_log = 30'b010101000100010011010000000100;
8'b00110100 : c0_log = 30'b010101000001000001100010010011;
8'b00110101 : c0_log = 30'b010100111101101001010001000110;
8'b00110110 : c0_log = 30'b010100111010010111100011010100;
8'b00110111 : c0_log = 30'b010100110111000101110101100011;
8'b00111000 : c0_log = 30'b010100110011110100000111110010;
8'b00111001 : c0_log = 30'b010100110000100010011010000000;
8'b00111010 : c0_log = 30'b010100101101010000101100001111;
8'b00111011 : c0_log = 30'b010100101001111110111110011101;
8'b00111100 : c0_log = 30'b010100100110110011110100000111;
8'b00111101 : c0_log = 30'b010100100011100010000110010110;
8'b00111110 : c0_log = 30'b010100100000010110111100000000;
8'b00111111 : c0_log = 30'b010100011101000101001110001110;
8'b01000000 : c0_log = 30'b010100011001111010000011111001;
8'b01000001 : c0_log = 30'b010100010110101110111001100011;
8'b01000010 : c0_log = 30'b010100010011100011101111001101;
8'b01000011 : c0_log = 30'b010100010000011000100100110111;
8'b01000100 : c0_log = 30'b010100001101001101011010100001;
8'b01000101 : c0_log = 30'b010100001010000010010000001011;
8'b01000110 : c0_log = 30'b010100000110110111000101110101;
8'b01000111 : c0_log = 30'b010100000011110010011110111011;
8'b01001000 : c0_log = 30'b010100000000100111010100100101;
8'b01001001 : c0_log = 30'b010011111101100010101101101010;
8'b01001010 : c0_log = 30'b010011111010011110000110110000;
8'b01001011 : c0_log = 30'b010011110111011001011111110110;
8'b01001100 : c0_log = 30'b010011110100001110010101100000;
8'b01001101 : c0_log = 30'b010011110001001001101110100101;
8'b01001110 : c0_log = 30'b010011101110000101000111101011;
8'b01001111 : c0_log = 30'b010011101011000111000100001100;
8'b01010000 : c0_log = 30'b010011101000000010011101010010;
8'b01010001 : c0_log = 30'b010011100100111101110110010111;
8'b01010010 : c0_log = 30'b010011100001111111110010111001;
8'b01010011 : c0_log = 30'b010011011110111011001011111110;
8'b01010100 : c0_log = 30'b010011011011111101001000011111;
8'b01010101 : c0_log = 30'b010011011000111000100001100101;
8'b01010110 : c0_log = 30'b010011010101111010011110000110;
8'b01010111 : c0_log = 30'b010011010010111100011010100111;
8'b01011000 : c0_log = 30'b010011001111111110010111001001;
8'b01011001 : c0_log = 30'b010011001101000000010011101010;
8'b01011010 : c0_log = 30'b010011001010000010010000001011;
8'b01011011 : c0_log = 30'b010011000111000100001100101100;
8'b01011100 : c0_log = 30'b010011000100000110001001001101;
8'b01011101 : c0_log = 30'b010011000001001110101001001010;
8'b01011110 : c0_log = 30'b010010111110010000100101101011;
8'b01011111 : c0_log = 30'b010010111011011001000101101000;
8'b01100000 : c0_log = 30'b010010111000011011000010001001;
8'b01100001 : c0_log = 30'b010010110101100011100010000110;
8'b01100010 : c0_log = 30'b010010110010101100000010000011;
8'b01100011 : c0_log = 30'b010010101111110100100001111111;
8'b01100100 : c0_log = 30'b010010101100110110011110100000;
8'b01100101 : c0_log = 30'b010010101001111110111110011101;
8'b01100110 : c0_log = 30'b010010100111000111011110011010;
8'b01100111 : c0_log = 30'b010010100100010110100001110010;
8'b01101000 : c0_log = 30'b010010100001011111000001101111;
8'b01101001 : c0_log = 30'b010010011110100111100001101100;
8'b01101010 : c0_log = 30'b010010011011110110100101000100;
8'b01101011 : c0_log = 30'b010010011000111111000101000001;
8'b01101100 : c0_log = 30'b010010010110001110001000011001;
8'b01101101 : c0_log = 30'b010010010011010110101000010110;
8'b01101110 : c0_log = 30'b010010010000100101101011101110;
8'b01101111 : c0_log = 30'b010010001101110100101111000110;
8'b01110000 : c0_log = 30'b010010001010111101001111000011;
8'b01110001 : c0_log = 30'b010010001000001100010010011011;
8'b01110010 : c0_log = 30'b010010000101011011010101110011;
8'b01110011 : c0_log = 30'b010010000010101010011001001100;
8'b01110100 : c0_log = 30'b010001111111111001011100100100;
8'b01110101 : c0_log = 30'b010001111101001111000011011000;
8'b01110110 : c0_log = 30'b010001111010011110000110110000;
8'b01110111 : c0_log = 30'b010001110111101101001010001000;
8'b01111000 : c0_log = 30'b010001110101000010110000111100;
8'b01111001 : c0_log = 30'b010001110010010001110100010100;
8'b01111010 : c0_log = 30'b010001101111100111011011001000;
8'b01111011 : c0_log = 30'b010001101100110110011110100000;
8'b01111100 : c0_log = 30'b010001101010001100000101010100;
8'b01111101 : c0_log = 30'b010001100111100001101100001000;
8'b01111110 : c0_log = 30'b010001100100110000101111100000;
8'b01111111 : c0_log = 30'b010001100010000110010110010100;
8'b10000000 : c0_log = 30'b010001011111011011111101001000;
8'b10000001 : c0_log = 30'b010001011100110001100011111100;
8'b10000010 : c0_log = 30'b010001011010000111001010110000;
8'b10000011 : c0_log = 30'b010001010111100011010100111111;
8'b10000100 : c0_log = 30'b010001010100111000111011110011;
8'b10000101 : c0_log = 30'b010001010010001110100010100111;
8'b10000110 : c0_log = 30'b010001001111101010101100110110;
8'b10000111 : c0_log = 30'b010001001101000000010011101010;
8'b10001000 : c0_log = 30'b010001001010010101111010011110;
8'b10001001 : c0_log = 30'b010001000111110010000100101101;
8'b10001010 : c0_log = 30'b010001000101001110001110111100;
8'b10001011 : c0_log = 30'b010001000010100011110101110000;
8'b10001100 : c0_log = 30'b010001                        ;
8'b10001101 : c0_log = 30'b010000111101011100001010001111;
8'b10001110 : c0_log = 30'b010000111010111000010100011110;
8'b10001111 : c0_log = 30'b010000111000010100011110101110;
8'b10010000 : c0_log = 30'b010000110101110000101000111101;
8'b10010001 : c0_log = 30'b010000110011001100110011001100;
8'b10010010 : c0_log = 30'b010000110000101000111101011100;
8'b10010011 : c0_log = 30'b010000101110000101000111101011;
8'b10010100 : c0_log = 30'b010000101011100001010001111010;
8'b10010101 : c0_log = 30'b010000101001000011111111100101;
8'b10010110 : c0_log = 30'b010000100110100000001001110101;
8'b10010111 : c0_log = 30'b010000100011111100010100000100;
8'b10011000 : c0_log = 30'b010000100001011111000001101111;
8'b10011001 : c0_log = 30'b010000011110111011001011111110;
8'b10011010 : c0_log = 30'b010000011100011101111001101001;
8'b10011011 : c0_log = 30'b010000011010000000100111010100;
8'b10011100 : c0_log = 30'b010000010111011100110001100011;
8'b10011101 : c0_log = 30'b010000010100111111011111001110;
8'b10011110 : c0_log = 30'b010000010010100010001100111001;
8'b10011111 : c0_log = 30'b010000010000000100111010100100;
8'b10100000 : c0_log = 30'b010000001101100111101000001111;
8'b10100001 : c0_log = 30'b010000001011001010010101111010;
8'b10100010 : c0_log = 30'b010000001000101101000011100101;
8'b10100011 : c0_log = 30'b010000000110001111110001010000;
8'b10100100 : c0_log = 30'b010000000011110010011110111011;
8'b10100101 : c0_log = 30'b010000000001011011110000000001;
8'b10100110 : c0_log = 30'b001111111110111101110011110000;
8'b10100111 : c0_log = 30'b001111111100100010011111010000;
8'b10101000 : c0_log = 30'b001111111010001000011110101000;
8'b10101001 : c0_log = 30'b001111110111101101110100000101;
8'b10101010 : c0_log = 30'b001111110101010100011101011010;
8'b10101011 : c0_log = 30'b001111110010111010011100110010;
8'b10101100 : c0_log = 30'b001111110000100001110000000100;
8'b10101101 : c0_log = 30'b001111101110001001000011010101;
8'b10101110 : c0_log = 30'b001111101011110000010110100111;
8'b10101111 : c0_log = 30'b001111101001011000010011110100;
8'b10110000 : c0_log = 30'b001111100111000000111010111110;
8'b10110001 : c0_log = 30'b001111100100101001100010001000;
8'b10110010 : c0_log = 30'b001111100010010010001001010011;
8'b10110011 : c0_log = 30'b001111011111111011011010011001;
8'b10110100 : c0_log = 30'b001111011101100101010101011100;
8'b10110101 : c0_log = 30'b001111011011001111010000011111;
8'b10110110 : c0_log = 30'b001111011000111001110101011110;
8'b10110111 : c0_log = 30'b001111010110100100011010011101;
8'b10111000 : c0_log = 30'b001111010100001111101001011000;
8'b10111001 : c0_log = 30'b001111010001111010111000010100;
8'b10111010 : c0_log = 30'b001111001111100110110001001100;
8'b10111011 : c0_log = 30'b001111001101010010101010000100;
8'b10111100 : c0_log = 30'b001111001010111111001100111000;
8'b10111101 : c0_log = 30'b001111001000101011101111101100;
8'b10111110 : c0_log = 30'b001111000110011000111100011101;
8'b10111111 : c0_log = 30'b001111000100000110001001001101;
8'b11000000 : c0_log = 30'b001111000001110011111111111010;
8'b11000001 : c0_log = 30'b001110111111100001110110100111;
8'b11000010 : c0_log = 30'b001110111101010000010111010000;
8'b11000011 : c0_log = 30'b001110111010111110110111111010;
8'b11000100 : c0_log = 30'b001110111000101110000010011111;
8'b11000101 : c0_log = 30'b001110110110011101001101000101;
8'b11000110 : c0_log = 30'b001110110100001101000001100111;
8'b11000111 : c0_log = 30'b001110110001111100110110001001;
8'b11001000 : c0_log = 30'b001110101111101101010100100111;
8'b11001001 : c0_log = 30'b001110101101011101110011000110;
8'b11001010 : c0_log = 30'b001110101011001110111011100000;
8'b11001011 : c0_log = 30'b001110101001000000000011111011;
8'b11001100 : c0_log = 30'b001110100110110001110110010010;
8'b11001101 : c0_log = 30'b001110100100100011101000101001;
8'b11001110 : c0_log = 30'b001110100010010101011011000000;
8'b11001111 : c0_log = 30'b001110100000000111110111010100;
8'b11010000 : c0_log = 30'b001110011101111010111101100100;
8'b11010001 : c0_log = 30'b001110011011101110000011110011;
8'b11010010 : c0_log = 30'b001110011001100001001010000011;
8'b11010011 : c0_log = 30'b001110010111010100111010001111;
8'b11010100 : c0_log = 30'b001110010101001000101010011011;
8'b11010101 : c0_log = 30'b001110010010111101000100100100;
8'b11010110 : c0_log = 30'b001110010000110001011110101100;
8'b11010111 : c0_log = 30'b001110001110100110100010110001;
8'b11011000 : c0_log = 30'b001110001100011011100110110110;
8'b11011001 : c0_log = 30'b001110001010010001010100110111;
8'b11011010 : c0_log = 30'b001110001000000111000010111000;
8'b11011011 : c0_log = 30'b001110000101111100110000111001;
8'b11011100 : c0_log = 30'b001110000011110011001000110111;
8'b11011101 : c0_log = 30'b001110000001101001100000110101;
8'b11011110 : c0_log = 30'b001101111111100000100010101110;
8'b11011111 : c0_log = 30'b001101111101010111100100101000;
8'b11100000 : c0_log = 30'b001101111011001111010000011111;
8'b11100001 : c0_log = 30'b001101111001000110111100010101;
8'b11100010 : c0_log = 30'b001101110110111111010010000111;
8'b11100011 : c0_log = 30'b001101110100110111100111111010;
8'b11100100 : c0_log = 30'b001101110010101111111101101101;
8'b11100101 : c0_log = 30'b001101110000101000111101011100;
8'b11100110 : c0_log = 30'b001101101110100001111101001011;
8'b11100111 : c0_log = 30'b001101101100011011100110110110;
8'b11101000 : c0_log = 30'b001101101010010101010000100001;
8'b11101001 : c0_log = 30'b001101101000001110111010001101;
8'b11101010 : c0_log = 30'b001101100110001001001101110100;
8'b11101011 : c0_log = 30'b001101100100000100001011011000;
8'b11101100 : c0_log = 30'b001101100001111110011111000000;
8'b11101101 : c0_log = 30'b001101011111111010000110100000;
8'b11101110 : c0_log = 30'b001101011101110101000100000100;
8'b11101111 : c0_log = 30'b001101011011110000101011100101;
8'b11110000 : c0_log = 30'b001101011001101100010011000101;
8'b11110001 : c0_log = 30'b001101010111101000100100100010;
8'b11110010 : c0_log = 30'b001101010101100100110101111111;
8'b11110011 : c0_log = 30'b001101010011100001110001011000;
8'b11110100 : c0_log = 30'b001101010001011110101100110001;
8'b11110101 : c0_log = 30'b001101001111011011101000001010;
8'b11110110 : c0_log = 30'b001101001101011001001101011111;
8'b11110111 : c0_log = 30'b001101001011010110110010110101;
8'b11111000 : c0_log = 30'b001101001001010101000010000111;
8'b11111001 : c0_log = 30'b001101000111010011010001011000;
8'b11111010 : c0_log = 30'b001101000101010001100000101010;
8'b11111011 : c0_log = 30'b001101000011010000011001111000;
8'b11111100 : c0_log = 30'b001101000001001111010011000110;
8'b11111101 : c0_log = 30'b001100111111001110110110010001;
8'b11111110 : c0_log = 30'b001100111101001110011001011011;
8'b11111111 : c0_log = 30'b001100111011001101111100100110;
endcase
end
endmodule
