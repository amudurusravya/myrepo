//------------------------------------------------------------------------------
// lookup table for cosine unit
// this will have c0,c1 stored and used for cosine coefficients lookup
// cosine_unit_lut.v
//
//------------------------------------------------------------------------------

module cosine_unit_lut(
  input [6:0] addr,
  output [11:0] c1_cosine_out,
  output [19:0] c0_cosine_out
);

reg [11:0] c1_cosine;
reg [19:0] c0_cosine;

assign c0_cosine_out = c0_cosine;
assign c1_cosine_out = c1_cosine;

always @(addr) begin
  case(addr)
7'b0000000 : c1_cosine = 12'b101111111111;
7'b0000001 : c1_cosine = 12'b110000000011;
7'b0000010 : c1_cosine = 12'b110000000110;
7'b0000011 : c1_cosine = 12'b110000001010;
7'b0000100 : c1_cosine = 12'b110000001101;
7'b0000101 : c1_cosine = 12'b110000010000;
7'b0000110 : c1_cosine = 12'b110000010011;
7'b0000111 : c1_cosine = 12'b110000010110;
7'b0001000 : c1_cosine = 12'b110000011001;
7'b0001001 : c1_cosine = 12'b110000011100;
7'b0001010 : c1_cosine = 12'b110000011111;
7'b0001011 : c1_cosine = 12'b110000100010;
7'b0001100 : c1_cosine = 12'b110000100101;
7'b0001101 : c1_cosine = 12'b110000101000;
7'b0001110 : c1_cosine = 12'b110000101011;
7'b0001111 : c1_cosine = 12'b110000101101;
7'b0010000 : c1_cosine = 12'b110000110000;
7'b0010001 : c1_cosine = 12'b110000110011;
7'b0010010 : c1_cosine = 12'b110000110101;
7'b0010011 : c1_cosine = 12'b110000111000;
7'b0010100 : c1_cosine = 12'b110000111010;
7'b0010101 : c1_cosine = 12'b110000111101;
7'b0010110 : c1_cosine = 12'b110000111111;
7'b0010111 : c1_cosine = 12'b110001000001;
7'b0011000 : c1_cosine = 12'b110001000100;
7'b0011001 : c1_cosine = 12'b110001000110;
7'b0011010 : c1_cosine = 12'b110001001000;
7'b0011011 : c1_cosine = 12'b110001001010;
7'b0011100 : c1_cosine = 12'b110001001100;
7'b0011101 : c1_cosine = 12'b110001001110;
7'b0011110 : c1_cosine = 12'b110001010000;
7'b0011111 : c1_cosine = 12'b110001010010;
7'b0100000 : c1_cosine = 12'b110001010100;
7'b0100001 : c1_cosine = 12'b110001010110;
7'b0100010 : c1_cosine = 12'b110001010111;
7'b0100011 : c1_cosine = 12'b110001011001;
7'b0100100 : c1_cosine = 12'b110001011011;
7'b0100101 : c1_cosine = 12'b110001011100;
7'b0100110 : c1_cosine = 12'b110001011110;
7'b0100111 : c1_cosine = 12'b110001011111;
7'b0101000 : c1_cosine = 12'b110001100000;
7'b0101001 : c1_cosine = 12'b110001100010;
7'b0101010 : c1_cosine = 12'b110001100011;
7'b0101011 : c1_cosine = 12'b110001100100;
7'b0101100 : c1_cosine = 12'b110001100101;
7'b0101101 : c1_cosine = 12'b110001100111;
7'b0101110 : c1_cosine = 12'b110001101000;
7'b0101111 : c1_cosine = 12'b110001101001;
7'b0110000 : c1_cosine = 12'b110001101001;
7'b0110001 : c1_cosine = 12'b110001101010;
7'b0110010 : c1_cosine = 12'b110001101011;
7'b0110011 : c1_cosine = 12'b110001101100;
7'b0110100 : c1_cosine = 12'b110001101101;
7'b0110101 : c1_cosine = 12'b110001101101;
7'b0110110 : c1_cosine = 12'b110001101110;
7'b0110111 : c1_cosine = 12'b110001101111;
7'b0111000 : c1_cosine = 12'b110001101111;
7'b0111001 : c1_cosine = 12'b110001101111;
7'b0111010 : c1_cosine = 12'b110001110000;
7'b0111011 : c1_cosine = 12'b110001110000;
7'b0111100 : c1_cosine = 12'b110001110000;
7'b0111101 : c1_cosine = 12'b110001110001;
7'b0111110 : c1_cosine = 12'b110001110001;
7'b0111111 : c1_cosine = 12'b110001110001;
7'b1000000 : c1_cosine = 12'b110001110001;
7'b1000001 : c1_cosine = 12'b110001110001;
7'b1000010 : c1_cosine = 12'b110001110001;
7'b1000011 : c1_cosine = 12'b110001110001;
7'b1000100 : c1_cosine = 12'b110001110000;
7'b1000101 : c1_cosine = 12'b110001110000;
7'b1000110 : c1_cosine = 12'b110001110000;
7'b1000111 : c1_cosine = 12'b110001101111;
7'b1001000 : c1_cosine = 12'b110001101111;
7'b1001001 : c1_cosine = 12'b110001101111;
7'b1001010 : c1_cosine = 12'b110001101110;
7'b1001011 : c1_cosine = 12'b110001101101;
7'b1001100 : c1_cosine = 12'b110001101101;
7'b1001101 : c1_cosine = 12'b110001101100;
7'b1001110 : c1_cosine = 12'b110001101011;
7'b1001111 : c1_cosine = 12'b110001101010;
7'b1010000 : c1_cosine = 12'b110001101001;
7'b1010001 : c1_cosine = 12'b110001101001;
7'b1010010 : c1_cosine = 12'b110001101000;
7'b1010011 : c1_cosine = 12'b110001100111;
7'b1010100 : c1_cosine = 12'b110001100101;
7'b1010101 : c1_cosine = 12'b110001100100;
7'b1010110 : c1_cosine = 12'b110001100011;
7'b1010111 : c1_cosine = 12'b110001100010;
7'b1011000 : c1_cosine = 12'b110001100000;
7'b1011001 : c1_cosine = 12'b110001011111;
7'b1011010 : c1_cosine = 12'b110001011110;
7'b1011011 : c1_cosine = 12'b110001011100;
7'b1011100 : c1_cosine = 12'b110001011011;
7'b1011101 : c1_cosine = 12'b110001011001;
7'b1011110 : c1_cosine = 12'b110001010111;
7'b1011111 : c1_cosine = 12'b110001010110;
7'b1100000 : c1_cosine = 12'b110001010100;
7'b1100001 : c1_cosine = 12'b110001010010;
7'b1100010 : c1_cosine = 12'b110001010000;
7'b1100011 : c1_cosine = 12'b110001001110;
7'b1100100 : c1_cosine = 12'b110001001100;
7'b1100101 : c1_cosine = 12'b110001001010;
7'b1100110 : c1_cosine = 12'b110001001000;
7'b1100111 : c1_cosine = 12'b110001000110;
7'b1101000 : c1_cosine = 12'b110001000100;
7'b1101001 : c1_cosine = 12'b110001000001;
7'b1101010 : c1_cosine = 12'b110000111111;
7'b1101011 : c1_cosine = 12'b110000111101;
7'b1101100 : c1_cosine = 12'b110000111010;
7'b1101101 : c1_cosine = 12'b110000111000;
7'b1101110 : c1_cosine = 12'b110000110101;
7'b1101111 : c1_cosine = 12'b110000110011;
7'b1110000 : c1_cosine = 12'b110000110000;
7'b1110001 : c1_cosine = 12'b110000101101;
7'b1110010 : c1_cosine = 12'b110000101011;
7'b1110011 : c1_cosine = 12'b110000101000;
7'b1110100 : c1_cosine = 12'b110000100101;
7'b1110101 : c1_cosine = 12'b110000100010;
7'b1110110 : c1_cosine = 12'b110000011111;
7'b1110111 : c1_cosine = 12'b110000011100;
7'b1111000 : c1_cosine = 12'b110000011001;
7'b1111001 : c1_cosine = 12'b110000010110;
7'b1111010 : c1_cosine = 12'b110000010011;
7'b1111011 : c1_cosine = 12'b110000010000;
7'b1111100 : c1_cosine = 12'b110000001101;
7'b1111101 : c1_cosine = 12'b110000001010;
7'b1111110 : c1_cosine = 12'b110000000110;
7'b1111111 : c1_cosine = 12'b110000000011;
endcase
end
always @(addr) begin
  case(addr)
7'b0000000 : c0_cosine = 20'b01000000000000000000;
7'b0000001 : c0_cosine = 20'b01000000011111111100;
7'b0000010 : c0_cosine = 20'b01000000111111000101;
7'b0000011 : c0_cosine = 20'b01000001011110001101;
7'b0000100 : c0_cosine = 20'b01000001111100111011;
7'b0000101 : c0_cosine = 20'b01000010011010110101;
7'b0000110 : c0_cosine = 20'b01000010111000101110;
7'b0000111 : c0_cosine = 20'b01000011010101110011;
7'b0001000 : c0_cosine = 20'b01000011110010111001;
7'b0001001 : c0_cosine = 20'b01000100001111001001;
7'b0001010 : c0_cosine = 20'b01000100101011000000;
7'b0001011 : c0_cosine = 20'b01000101000110110111;
7'b0001100 : c0_cosine = 20'b01000101100001111001;
7'b0001101 : c0_cosine = 20'b01000101111100100001;
7'b0001110 : c0_cosine = 20'b01000110010110101110;
7'b0001111 : c0_cosine = 20'b01000110110000100010;
7'b0010000 : c0_cosine = 20'b01000111001001100001;
7'b0010001 : c0_cosine = 20'b01000111100010100000;
7'b0010010 : c0_cosine = 20'b01000111111010101011;
7'b0010011 : c0_cosine = 20'b01001000010010110101;
7'b0010100 : c0_cosine = 20'b01001000101010001100;
7'b0010101 : c0_cosine = 20'b01001001000001001000;
7'b0010110 : c0_cosine = 20'b01001001010111001111;
7'b0010111 : c0_cosine = 20'b01001001101101010111;
7'b0011000 : c0_cosine = 20'b01001010000010101010;
7'b0011001 : c0_cosine = 20'b01001010010111100011;
7'b0011010 : c0_cosine = 20'b01001010101100000010;
7'b0011011 : c0_cosine = 20'b01001011000000000110;
7'b0011100 : c0_cosine = 20'b01001011010011110000;
7'b0011101 : c0_cosine = 20'b01001011100110100110;
7'b0011110 : c0_cosine = 20'b01001011111001000010;
7'b0011111 : c0_cosine = 20'b01001100001011000011;
7'b0100000 : c0_cosine = 20'b01001100011100101011;
7'b0100001 : c0_cosine = 20'b01001100101101011101;
7'b0100010 : c0_cosine = 20'b01001100111101110110;
7'b0100011 : c0_cosine = 20'b01001101001101110100;
7'b0100100 : c0_cosine = 20'b01001101011101011000;
7'b0100101 : c0_cosine = 20'b01001101101100001000;
7'b0100110 : c0_cosine = 20'b01001101111010011110;
7'b0100111 : c0_cosine = 20'b01001110001000011001;
7'b0101000 : c0_cosine = 20'b01001110010101100000;
7'b0101001 : c0_cosine = 20'b01001110100010001100;
7'b0101010 : c0_cosine = 20'b01001110101110011111;
7'b0101011 : c0_cosine = 20'b01001110111010010111;
7'b0101100 : c0_cosine = 20'b01001111000101011011;
7'b0101101 : c0_cosine = 20'b01001111010000000100;
7'b0101110 : c0_cosine = 20'b01001111011010010100;
7'b0101111 : c0_cosine = 20'b01001111100011101111;
7'b0110000 : c0_cosine = 20'b01001111101100101111;
7'b0110001 : c0_cosine = 20'b01001111110101010110;
7'b0110010 : c0_cosine = 20'b01001111111101001000;
7'b0110011 : c0_cosine = 20'b01010000000100100000;
7'b0110100 : c0_cosine = 20'b01010000001011011110;
7'b0110101 : c0_cosine = 20'b01010000010001100111;
7'b0110110 : c0_cosine = 20'b01010000010111010110;
7'b0110111 : c0_cosine = 20'b01010000011100101011;
7'b0111000 : c0_cosine = 20'b01010000100001001011;
7'b0111001 : c0_cosine = 20'b01010000100101101011;
7'b0111010 : c0_cosine = 20'b01010000101000111101;
7'b0111011 : c0_cosine = 20'b01010000101100001111;
7'b0111100 : c0_cosine = 20'b01010000101110101100;
7'b0111101 : c0_cosine = 20'b01010000110000010101;
7'b0111110 : c0_cosine = 20'b01010000110001111110;
7'b0111111 : c0_cosine = 20'b01010000110010110010;
7'b1000000 : c0_cosine = 20'b01010000110010110010;
7'b1000001 : c0_cosine = 20'b01010000110010110010;
7'b1000010 : c0_cosine = 20'b01010000110001111110;
7'b1000011 : c0_cosine = 20'b01010000110000010101;
7'b1000100 : c0_cosine = 20'b01010000101110101100;
7'b1000101 : c0_cosine = 20'b01010000101100001111;
7'b1000110 : c0_cosine = 20'b01010000101000111101;
7'b1000111 : c0_cosine = 20'b01010000100101010001;
7'b1001000 : c0_cosine = 20'b01010000100001001011;
7'b1001001 : c0_cosine = 20'b01010000011100101011;
7'b1001010 : c0_cosine = 20'b01010000010111010110;
7'b1001011 : c0_cosine = 20'b01010000010001100111;
7'b1001100 : c0_cosine = 20'b01010000001011011110;
7'b1001101 : c0_cosine = 20'b01010000000100100000;
7'b1001110 : c0_cosine = 20'b01001111111101001000;
7'b1001111 : c0_cosine = 20'b01001111110101010110;
7'b1010000 : c0_cosine = 20'b01001111101100101111;
7'b1010001 : c0_cosine = 20'b01001111100011101111;
7'b1010010 : c0_cosine = 20'b01001111011001111010;
7'b1010011 : c0_cosine = 20'b01001111010000000100;
7'b1010100 : c0_cosine = 20'b01001111000101011011;
7'b1010101 : c0_cosine = 20'b01001110111010010111;
7'b1010110 : c0_cosine = 20'b01001110101110011111;
7'b1010111 : c0_cosine = 20'b01001110100010001100;
7'b1011000 : c0_cosine = 20'b01001110010101100000;
7'b1011001 : c0_cosine = 20'b01001110000111111111;
7'b1011010 : c0_cosine = 20'b01001101111010011110;
7'b1011011 : c0_cosine = 20'b01001101101100001000;
7'b1011100 : c0_cosine = 20'b01001101011100111110;
7'b1011101 : c0_cosine = 20'b01001101001101110100;
7'b1011110 : c0_cosine = 20'b01001100111101110110;
7'b1011111 : c0_cosine = 20'b01001100101101011101;
7'b1100000 : c0_cosine = 20'b01001100011100010000;
7'b1100001 : c0_cosine = 20'b01001100001011000011;
7'b1100010 : c0_cosine = 20'b01001011111001000010;
7'b1100011 : c0_cosine = 20'b01001011100110100110;
7'b1100100 : c0_cosine = 20'b01001011010011010110;
7'b1100101 : c0_cosine = 20'b01001011000000000110;
7'b1100110 : c0_cosine = 20'b01001010101100000010;
7'b1100111 : c0_cosine = 20'b01001010010111100011;
7'b1101000 : c0_cosine = 20'b01001010000010101010;
7'b1101001 : c0_cosine = 20'b01001001101100111101;
7'b1101010 : c0_cosine = 20'b01001001010111001111;
7'b1101011 : c0_cosine = 20'b01001001000000101101;
7'b1101100 : c0_cosine = 20'b01001000101001110001;
7'b1101101 : c0_cosine = 20'b01001000010010011011;
7'b1101110 : c0_cosine = 20'b01000111111010101011;
7'b1101111 : c0_cosine = 20'b01000111100010000110;
7'b1110000 : c0_cosine = 20'b01000111001001100001;
7'b1110001 : c0_cosine = 20'b01000110110000001000;
7'b1110010 : c0_cosine = 20'b01000110010110010100;
7'b1110011 : c0_cosine = 20'b01000101111100000110;
7'b1110100 : c0_cosine = 20'b01000101100001011111;
7'b1110101 : c0_cosine = 20'b01000101000110011100;
7'b1110110 : c0_cosine = 20'b01000100101011000000;
7'b1110111 : c0_cosine = 20'b01000100001111001001;
7'b1111000 : c0_cosine = 20'b01000011110010011110;
7'b1111001 : c0_cosine = 20'b01000011010101110011;
7'b1111010 : c0_cosine = 20'b01000010111000010100;
7'b1111011 : c0_cosine = 20'b01000010011010110101;
7'b1111100 : c0_cosine = 20'b01000001111100100001;
7'b1111101 : c0_cosine = 20'b01000001011101110011;
7'b1111110 : c0_cosine = 20'b01000000111111000101;
7'b1111111 : c0_cosine = 20'b01000000011111100010;
endcase
end
endmodule
